module RISC_V(
  input clk, reset_n
);
endmodule
